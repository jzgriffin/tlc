(* TLC in Coq
 *
 * Module: tlc.utility.all_utility
 * Purpose: Exports the entire utility module by exporting all submodules.
 *
 * The utility module contains types and functions that are not part of TLC
 * but are used in its implementation.  Each submodule typically contains a
 * single type, for which it is named, or a set of functions defined for a
 * particular existing type.  For example, the seq submodule contains
 * functions augmenting the ssreflect seq type, while the result type defines
 * the result monad type.
 *
 * Included in this module is the functor -> applicative functor -> monad
 * hierarchy of typeclasses that appears in Haskell.
 *)

Require Export tlc.utility.applicative.
Require Export tlc.utility.ascii.
Require Export tlc.utility.functor.
Require Export tlc.utility.monad.
Require Export tlc.utility.option.
Require Export tlc.utility.partial_map.
Require Export tlc.utility.result.
Require Export tlc.utility.seq.
Require Export tlc.utility.set.
Require Export tlc.utility.string.
